//-------------------------------------------------------------------------
//      lab8.sv                                                          --
//      Christine Chen                                                   --
//      Fall 2014                                                        --
//                                                                       --
//      Modified by Po-Han Huang                                         --
//      10/06/2017                                                       --
//                                                                       --
//      Fall 2017 Distribution                                           --
//                                                                       --
//      For use with ECE 385 Lab 8                                       --
//      UIUC ECE Department                                              --
//-------------------------------------------------------------------------


module lab8( input               CLOCK_50,
             input        [3:0]  KEY,          //bit 0 is set up as Reset
             output logic [6:0]  HEX0, HEX1,
				 output logic [3:0]  LEDG,				//added
             // VGA Interface
             output logic [7:0]  VGA_R,        //VGA Red
                                 VGA_G,        //VGA Green
                                 VGA_B,        //VGA Blue
             output logic        VGA_CLK,      //VGA Clock
                                 VGA_SYNC_N,   //VGA Sync signal
                                 VGA_BLANK_N,  //VGA Blank signal
                                 VGA_VS,       //VGA virtical sync signal
                                 VGA_HS,       //VGA horizontal sync signal
             // CY7C67200 Interface
             inout  wire  [15:0] OTG_DATA,     //CY7C67200 Data bus 16 Bits
             output logic [1:0]  OTG_ADDR,     //CY7C67200 Address 2 Bits
             output logic        OTG_CS_N,     //CY7C67200 Chip Select
                                 OTG_RD_N,     //CY7C67200 Write
                                 OTG_WR_N,     //CY7C67200 Read
                                 OTG_RST_N,    //CY7C67200 Reset
             input               OTG_INT,      //CY7C67200 Interrupt
             // SDRAM Interface for Nios II Software
             output logic [12:0] DRAM_ADDR,    //SDRAM Address 13 Bits
             inout  wire  [31:0] DRAM_DQ,      //SDRAM Data 32 Bits
             output logic [1:0]  DRAM_BA,      //SDRAM Bank Address 2 Bits
             output logic [3:0]  DRAM_DQM,     //SDRAM Data Mast 4 Bits
             output logic        DRAM_RAS_N,   //SDRAM Row Address Strobe
                                 DRAM_CAS_N,   //SDRAM Column Address Strobe
                                 DRAM_CKE,     //SDRAM Clock Enable
                                 DRAM_WE_N,    //SDRAM Write Enable
                                 DRAM_CS_N,    //SDRAM Chip Select
                                 DRAM_CLK      //SDRAM Clock
                    );

    logic Reset_h, Clk, Run_h;
    logic [7:0] keycode;

	 //added variables
    logic [9:0] Draw_X, Draw_Y;
	 logic is_ball;
	 logic [3:0] LEDA;

    assign Clk = CLOCK_50;
    always_ff @ (posedge Clk) begin
        Reset_h <= ~(KEY[0]);        // The push buttons are active low
		  Run_h <= ~(KEY[1]);
	end

    logic [1:0] hpi_addr;
    logic [15:0] hpi_data_in, hpi_data_out;
    logic hpi_r, hpi_w, hpi_cs, hpi_reset;


	 assign LEDG = LEDA;

    // Interface between NIOS II and EZ-OTG chip
    hpi_io_intf hpi_io_inst(
                            .Clk(Clk),
                            .Reset(Reset_h),
                            // signals connected to NIOS II
                            .from_sw_address(hpi_addr),
                            .from_sw_data_in(hpi_data_in),
                            .from_sw_data_out(hpi_data_out),
                            .from_sw_r(hpi_r),
                            .from_sw_w(hpi_w),
                            .from_sw_cs(hpi_cs),
                            .from_sw_reset(hpi_reset),
                            // signals connected to EZ-OTG chip
                            .OTG_DATA(OTG_DATA),
                            .OTG_ADDR(OTG_ADDR),
                            .OTG_RD_N(OTG_RD_N),
                            .OTG_WR_N(OTG_WR_N),
                            .OTG_CS_N(OTG_CS_N),
                            .OTG_RST_N(OTG_RST_N)
    );

     // You need to make sure that the port names here match the ports in Qsys-generated codes.
     lab8_soc nios_system(
                             .clk_clk(Clk),
                             .reset_reset_n(1'b1),    // Never reset NIOS
                             .sdram_wire_addr(DRAM_ADDR),
                             .sdram_wire_ba(DRAM_BA),
                             .sdram_wire_cas_n(DRAM_CAS_N),
                             .sdram_wire_cke(DRAM_CKE),
                             .sdram_wire_cs_n(DRAM_CS_N),
                             .sdram_wire_dq(DRAM_DQ),
                             .sdram_wire_dqm(DRAM_DQM),
                             .sdram_wire_ras_n(DRAM_RAS_N),
                             .sdram_wire_we_n(DRAM_WE_N),
                             .sdram_clk_clk(DRAM_CLK),
                             .keycode_export(keycode),
                             .otg_hpi_address_export(hpi_addr),
                             .otg_hpi_data_in_port(hpi_data_in),
                             .otg_hpi_data_out_port(hpi_data_out),
                             .otg_hpi_cs_export(hpi_cs),
                             .otg_hpi_r_export(hpi_r),
                             .otg_hpi_w_export(hpi_w),
                             .otg_hpi_reset_export(hpi_reset)
    );

    // Use PLL to generate the 25MHZ VGA_CLK.
    // You will have to generate it on your own in simulation.
    vga_clk vga_clk_instance(.inclk0(Clk), .c0(VGA_CLK));

    // TODO: Fill in the connections for the rest of the modules
    VGA_controller vga_controller_instance(.Clk(Clk),
														.Reset(Reset_h),
														.VGA_HS(VGA_HS),
														.VGA_VS(VGA_VS),
														.VGA_CLK(VGA_CLK),
														.VGA_BLANK_N(VGA_BLANK_N),
														.VGA_SYNC_N(VGA_SYNC_N),
														.DrawX(Draw_X),
														.DrawY(Draw_Y));

	always_comb
	begin
	LEDA = 4'b0000;

	case (keycode)

	8'h001A: LEDA = 4'b1000; // up 1A
	8'h0016: LEDA = 4'b0001; // down 0016
	8'h0004: LEDA = 4'b0100; // left 0004
	8'h0007: LEDA = 4'b0010; // right 0007
	default: LEDA = 4'b0000;

	endcase
	end

    // Which signal should be frame_clk?  VGA CLK? VGA_VS Instead.
   ball ball_instance( .Clk(Clk),
	                    .Reset(Reset_h),
							  .Run(Run_h),
	                    .frame_clk(VGA_VS),
							  //.blank(VGA_BLANK_N),
							  .go(playerSig),
	                    .DrawX(Draw_X),
							  .DrawY(Draw_Y),
							  .xcent(10'd498),
							  .ycent(10'd418),
							  .button(delaypress),
	                    .is_ball(is_boll),
							  .turndone(playerdone)
	);

	logic is_mummy, is_boll;

	mummy mum_instance( .Clk(Clk),
	                    .Reset(Reset_h),
							  .Run(Run_h),
	                    .frame_clk(VGA_VS),
							  //.blank(VGA_BLANK_N),
							  .go(mummySig),
							  .go2(mummySig2),
	                    .DrawX(Draw_X),
							  .DrawY(Draw_Y),
							  .xcent(10'd141),
							  .ycent(10'd61),
							  .button(delaypress),
	                    .is_ball(is_mummy),
							  .turn1done(mummydone1),
							  .turn2done(mummydone2)
	);



   color_mapper color_instance( .is_ball(is_boll),
										  .is_mum(is_mummy),
										  .DrawX(Draw_X),
										  .DrawY(Draw_Y),
										  .VGA_R(VGA_R),
										  .VGA_G(VGA_G),
										  .VGA_B(VGA_B)
	 );

logic playerSig, mummySig, mummySig2, playerdone, mummydone1, mummydone2;

logic begincounting, donecounting, delaypress;

module timer(.Clk(Clk), .Reset(Reset_h), .enable(begincounting), .keyin(LEDG), .keyout(delaypress),
              .ticktock(donecounting));

FSM finite (
.Clk(Clk),
.Reset(Reset_h),
.Run(Run_h),


.playdon(playerdone), .mumdon1(mummydone1), .mumdon2(mummydone2), .VS(VGA_VS), //Tell the FSM the player has finished inputing a move //Tell the FSM the enemy has made a move
// 1 is enemy turn, 0 is player turn

//input logic win,
//input logic loss,
//input logic cont,

.playerSignal(playerSig),
.mummySignal(mummySig), .mummySignal2(mummySig2),
.startcounting(begincounting), .delayachieved(donecounting)


//output logic opening,
//output logic gameover, //output signals to stop the game
//output logic winner



);

    // Display keycode on hex display
    HexDriver hex_inst_0 (keycode[3:0], HEX0);
    HexDriver hex_inst_1 (keycode[7:4], HEX1);

    /**************************************************************************************
        ATTENTION! Please answer the following quesiton in your lab report! Points will be allocated for the answers!
        Hidden Question #1/2:
        What are the advantages and/or disadvantages of using a USB interface over PS/2 interface to
             connect to the keyboard? List any two.  Give an answer in your Post-Lab.
    **************************************************************************************/
endmodule






////-------------------------------------------------------------------------
////      lab8.sv                                                          --
////      Christine Chen                                                   --
////      Fall 2014                                                        --
////                                                                       --
////      Modified by Po-Han Huang                                         --
////      10/06/2017                                                       --
////                                                                       --
////      Fall 2017 Distribution                                           --
////                                                                       --
////      For use with ECE 385 Lab 8                                       --
////      UIUC ECE Department                                              --
////-------------------------------------------------------------------------
//
//
//module lab8( input               CLOCK_50,
//             input        [3:0]  KEY,          //bit 0 is set up as Reset
//             output logic [6:0]  HEX0, HEX1,
//				 output logic [3:0]  LEDG,				//added
//             // VGA Interface
//             output logic [7:0]  VGA_R,        //VGA Red
//                                 VGA_G,        //VGA Green
//                                 VGA_B,        //VGA Blue
//             output logic        VGA_CLK,      //VGA Clock
//                                 VGA_SYNC_N,   //VGA Sync signal
//                                 VGA_BLANK_N,  //VGA Blank signal
//                                 VGA_VS,       //VGA virtical sync signal
//                                 VGA_HS,       //VGA horizontal sync signal
//             // CY7C67200 Interface
//             inout  wire  [15:0] OTG_DATA,     //CY7C67200 Data bus 16 Bits
//             output logic [1:0]  OTG_ADDR,     //CY7C67200 Address 2 Bits
//             output logic        OTG_CS_N,     //CY7C67200 Chip Select
//                                 OTG_RD_N,     //CY7C67200 Write
//                                 OTG_WR_N,     //CY7C67200 Read
//                                 OTG_RST_N,    //CY7C67200 Reset
//             input               OTG_INT,      //CY7C67200 Interrupt
//             // SDRAM Interface for Nios II Software
//             output logic [12:0] DRAM_ADDR,    //SDRAM Address 13 Bits
//             inout  wire  [31:0] DRAM_DQ,      //SDRAM Data 32 Bits
//             output logic [1:0]  DRAM_BA,      //SDRAM Bank Address 2 Bits
//             output logic [3:0]  DRAM_DQM,     //SDRAM Data Mast 4 Bits
//             output logic        DRAM_RAS_N,   //SDRAM Row Address Strobe
//                                 DRAM_CAS_N,   //SDRAM Column Address Strobe
//                                 DRAM_CKE,     //SDRAM Clock Enable
//                                 DRAM_WE_N,    //SDRAM Write Enable
//                                 DRAM_CS_N,    //SDRAM Chip Select
//                                 DRAM_CLK      //SDRAM Clock
//                    );
//
//    logic Reset_h, Clk;
//    logic [7:0] keycode;
//
//	 //added variables
//    logic [9:0] Draw_X, Draw_Y;
//	 logic is_ball;
//	 logic [3:0] LEDA;
//
//    assign Clk = CLOCK_50;
//    always_ff @ (posedge Clk) begin
//        Reset_h <= ~(KEY[0]);        // The push buttons are active low
//    end
//
//    logic [1:0] hpi_addr;
//    logic [15:0] hpi_data_in, hpi_data_out;
//    logic hpi_r, hpi_w, hpi_cs, hpi_reset;
//
//
//	 assign LEDG = LEDA;
//
//    // Interface between NIOS II and EZ-OTG chip
//    hpi_io_intf hpi_io_inst(
//                            .Clk(Clk),
//                            .Reset(Reset_h),
//                            // signals connected to NIOS II
//                            .from_sw_address(hpi_addr),
//                            .from_sw_data_in(hpi_data_in),
//                            .from_sw_data_out(hpi_data_out),
//                            .from_sw_r(hpi_r),
//                            .from_sw_w(hpi_w),
//                            .from_sw_cs(hpi_cs),
//                            .from_sw_reset(hpi_reset),
//                            // signals connected to EZ-OTG chip
//                            .OTG_DATA(OTG_DATA),
//                            .OTG_ADDR(OTG_ADDR),
//                            .OTG_RD_N(OTG_RD_N),
//                            .OTG_WR_N(OTG_WR_N),
//                            .OTG_CS_N(OTG_CS_N),
//                            .OTG_RST_N(OTG_RST_N)
//    );
//
//     // You need to make sure that the port names here match the ports in Qsys-generated codes.
//     lab8_soc nios_system(
//                             .clk_clk(Clk),
//                             .reset_reset_n(1'b1),    // Never reset NIOS
//                             .sdram_wire_addr(DRAM_ADDR),
//                             .sdram_wire_ba(DRAM_BA),
//                             .sdram_wire_cas_n(DRAM_CAS_N),
//                             .sdram_wire_cke(DRAM_CKE),
//                             .sdram_wire_cs_n(DRAM_CS_N),
//                             .sdram_wire_dq(DRAM_DQ),
//                             .sdram_wire_dqm(DRAM_DQM),
//                             .sdram_wire_ras_n(DRAM_RAS_N),
//                             .sdram_wire_we_n(DRAM_WE_N),
//                             .sdram_clk_clk(DRAM_CLK),
//                             .keycode_export(keycode),
//                             .otg_hpi_address_export(hpi_addr),
//                             .otg_hpi_data_in_port(hpi_data_in),
//                             .otg_hpi_data_out_port(hpi_data_out),
//                             .otg_hpi_cs_export(hpi_cs),
//                             .otg_hpi_r_export(hpi_r),
//                             .otg_hpi_w_export(hpi_w),
//                             .otg_hpi_reset_export(hpi_reset)
//    );
//
//    // Use PLL to generate the 25MHZ VGA_CLK.
//    // You will have to generate it on your own in simulation.
//    vga_clk vga_clk_instance(.inclk0(Clk), .c0(VGA_CLK));
//
//    // TODO: Fill in the connections for the rest of the modules
//    VGA_controller vga_controller_instance(.Clk(Clk),
//														.Reset(Reset_h),
//														.VGA_HS(VGA_HS),
//														.VGA_VS(VGA_VS),
//														.VGA_CLK(VGA_CLK),
//														.VGA_BLANK_N(VGA_BLANK_N),
//														.VGA_SYNC_N(VGA_SYNC_N),
//														.DrawX(Draw_X),
//														.DrawY(Draw_Y));
//
//	always_comb
//	begin
//	LEDA = 4'b0000;
//
//	case (keycode)
//
//	8'h001A: LEDA = 4'b1000; // up 1A
//	8'h0016: LEDA = 4'b0001; // down 0016
//	8'h0004: LEDA = 4'b0100; // left 0004
//	8'h0007: LEDA = 4'b0010; // right 0007
//	default: LEDA = 4'b0000;
//
//	endcase
//	end
//
//
//    // Which signal should be frame_clk?  VGA CLK? VGA_VS Instead.
//   ball ball_instance( .Clk(Clk),
//	                    .Reset(Reset_h),
//	                    .frame_clk(VGA_VS),
//	                    .DrawX(Draw_X),
//							  .DrawY(Draw_Y),
//							  .button(LEDG),
//	                    .is_ball(is_ball)
//	);
//
//
//   color_mapper color_instance( .is_ball(is_ball),
//										  .DrawX(Draw_X),
//										  .DrawY(Draw_Y),
//										  .VGA_R(VGA_R),
//										  .VGA_G(VGA_G),
//										  .VGA_B(VGA_B)
//	 );
//
//    // Display keycode on hex display
//    HexDriver hex_inst_0 (keycode[3:0], HEX0);
//    HexDriver hex_inst_1 (keycode[7:4], HEX1);
//
//    /**************************************************************************************
//        ATTENTION! Please answer the following quesiton in your lab report! Points will be allocated for the answers!
//        Hidden Question #1/2:
//        What are the advantages and/or disadvantages of using a USB interface over PS/2 interface to
//             connect to the keyboard? List any two.  Give an answer in your Post-Lab.
//    **************************************************************************************/
//endmodule
